-- very simple tb to create an inboud and an outbound transactions.

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
USE ieee.numeric_std.ALL; 

entity tb is
end tb;

architecture tb of tb is
    -- change here if you want to send more packets
    constant N_PACKETS : integer := 4; 
    -- change here if you want to send longer packets
    constant MAX_FLITS : integer := 3;

	signal clock:    std_logic := '0';
	signal reset:    std_logic;  

	-- slave local port
    signal validL_i : std_logic;
    signal dataL_i  : std_logic_vector(31 downto 0);
    signal readyL_o : std_logic;                    

	-- master local port
    signal validL_o : std_logic;                    
    signal dataL_o  : std_logic_vector(31 downto 0);
    signal readyL_i : std_logic;                    
    signal lastL_o  : std_logic;                    
	
    -- other master ports
    signal validE_o : std_logic;                    
    signal dataE_o  : std_logic_vector(31 downto 0);
    signal readyE_i : std_logic;                    
    signal lastE_o  : std_logic;                    
            
    signal validW_o : std_logic;                    
    signal dataW_o  : std_logic_vector(31 downto 0);
    signal readyW_i : std_logic;                    
    signal lastW_o  : std_logic;                    
            
    signal validN_o : std_logic;                    
    signal dataN_o  : std_logic_vector(31 downto 0);
    signal readyN_i : std_logic;                    
    signal lastN_o  : std_logic;                    
            
    signal validS_o : std_logic;                    
    signal dataS_o  : std_logic_vector(31 downto 0);
    signal readyS_i : std_logic;                    
    signal lastS_o  : std_logic;                    
            
	
	
	
	-- send one work according to the AXI Streaming master protocol
	procedure SendFlit(signal clock  : in  std_logic;
	                   constant flit : in  std_logic_vector(31 downto 0);
	                   --- AXI master streaming 
	                   signal data   : out std_logic_vector(31 downto 0);
	                   signal valid  : out std_logic;
	                   signal ready  : in  std_logic
	                   ) is
	begin
		wait until rising_edge(clock);
		-- If both the AXI interface and the router runs at the rising edge, then it is necessary to add 
		--   a delay at the inputs. The solution was to put an inverted in the clock in the Router_Board entity. 
		-- This way the delay is not necessary and it is also not necessary to change the router's vhdl   
        data <= flit;
        valid <= '1';
        wait for 8ns; -- simulate delay at the primary inputs
        while ready /= '1' loop
             wait until falling_edge(clock); -- data is buffered at the falling edge
        end loop;	
	end procedure;
	
	
begin

	reset <= '1', '0' after 100 ns; -- active low

    -- 50 MHz, as the default freq generated by the PS
	process
	begin
		clock <= not clock;
		wait for 10 ns;
		clock <= not clock;
		wait for 10 ns;
	end process;
	
	-- master ports are always ready to receive
	readyE_i <= '1';
	readyN_i <= '1';
	readyW_i <= '1';
	readyS_i <= '1';
	readyL_i <= '1';

    ----------------------------------------------------
    -- testing the flow from the slave port to the Sink LEDs
    ----------------------------------------------------
    process
        -- it sends N_PACKETS packets of max size of of MAX_FLITS 
        type packet_vet_t is array (0 to N_PACKETS-1, 0 to MAX_FLITS+1) of std_logic_vector(31 downto 0);
        constant packet_vet : packet_vet_t := 
            (
                (x"00000201", x"00000001", x"00001234", x"00000000", x"00000000"), -- send it to the east
                (x"00000102", x"00000001", x"00004321", x"00000000", x"00000000"), -- send it to the north
                (x"00000001", x"00000003", x"11111111", x"22222222", x"33333333"), -- send it to the west
                (x"00000100", x"00000003", x"44444444", x"55555555", x"66666666")  -- send it to the south
            );
         variable num_flits : integer;
	begin
		validL_i <= '0';
		dataL_i <= (others => '0');
		wait for 200 ns;
		wait until rising_edge(clock);
		
		for p in 0 to N_PACKETS-1 loop
		  -- send header
		  SendFlit(clock,packet_vet(p,0),dataL_i,validL_i,readyL_o);
		  -- send size
		  SendFlit(clock,packet_vet(p,1),dataL_i,validL_i,readyL_o);
		  num_flits := to_integer(signed(packet_vet(p,1))) ;
		  -- send payload
		  for f in 2 to num_flits+1 loop
		      SendFlit(clock,packet_vet(p,f),dataL_i,validL_i,readyL_o);
		  end loop;
		-- end of the packet transfer
          wait until rising_edge(clock);
          wait for 4 ns;
          validL_i <= '0';
          dataL_i <= (others => '0');
          -- wait a while to start the next packet transfer 
          wait for 100 ns;
		end loop;
		
		-- blobk here. do not send it again
		wait;
	end process;


 router: entity work.RouterCC
  port map ( 
        clock    => clock,
        reset    => reset,
        -- AXI slave streaming interfaces
        validE_i => '0',
        dataE_i  => (others => '0'),
        readyE_o => open,          

        validW_i => '0',           
        dataW_i  => (others => '0'),
        readyW_o => open,          

        validN_i => '0',           
        dataN_i  => (others => '0'),
        readyN_o => open,          

        validS_i => '0',           
        dataS_i  => (others => '0'),
        readyS_o => open,          

        validL_i => validL_i,
        dataL_i  => dataL_i ,
        readyL_o => readyL_o,

        -- AXI master streaming interfaces
        validE_o => validE_o,
        dataE_o  => dataE_o ,
        readyE_i => readyE_i,
        lastE_o  => lastE_o ,

        validW_o => validW_o,
        dataW_o  => dataW_o ,
        readyW_i => readyW_i,
        lastW_o  => lastW_o ,

        validN_o => validN_o,
        dataN_o  => dataN_o ,
        readyN_i => readyN_i,
        lastN_o  => lastN_o ,

        validS_o => validS_o,
        dataS_o  => dataS_o ,
        readyS_i => readyS_i,
        lastS_o  => lastS_o ,

        validL_o => validL_o,
        dataL_o  => dataL_o ,
        readyL_i => readyL_i,
        lastL_o  => lastL_o 
	);
	
end tb;

